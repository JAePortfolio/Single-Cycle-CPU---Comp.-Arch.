library verilog;
use verilog.vl_types.all;
entity Arena_bitwiseor_vlg_vec_tst is
end Arena_bitwiseor_vlg_vec_tst;

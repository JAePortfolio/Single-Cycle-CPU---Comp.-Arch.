library verilog;
use verilog.vl_types.all;
entity Arena_Shift_Left_32bit_vlg_vec_tst is
end Arena_Shift_Left_32bit_vlg_vec_tst;

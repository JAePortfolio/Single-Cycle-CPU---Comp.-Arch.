library verilog;
use verilog.vl_types.all;
entity Arena_muxLPM_vlg_check_tst is
    port(
        Arena_result    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_muxLPM_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_fullAdder_vlg_vec_tst is
end Arena_fullAdder_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_ALU_Control_VHDL_vlg_vec_tst is
end Arena_ALU_Control_VHDL_vlg_vec_tst;

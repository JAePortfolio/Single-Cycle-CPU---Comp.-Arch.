library verilog;
use verilog.vl_types.all;
entity Arena_DataMemory_vlg_vec_tst is
end Arena_DataMemory_vlg_vec_tst;

-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: Arena_parallelAdder.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Arena_parallelAdder IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
	);
END Arena_parallelAdder;


ARCHITECTURE SYN OF arena_paralleladder IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire2	: ALTERA_MF_LOGIC_2D (16 DOWNTO 0, 0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (0 DOWNTO 0);

BEGIN
	sub_wire18    <= data0x(0 DOWNTO 0);
	sub_wire17    <= data1x(0 DOWNTO 0);
	sub_wire16    <= data2x(0 DOWNTO 0);
	sub_wire15    <= data3x(0 DOWNTO 0);
	sub_wire14    <= data4x(0 DOWNTO 0);
	sub_wire13    <= data5x(0 DOWNTO 0);
	sub_wire12    <= data6x(0 DOWNTO 0);
	sub_wire11    <= data7x(0 DOWNTO 0);
	sub_wire10    <= data8x(0 DOWNTO 0);
	sub_wire9    <= data9x(0 DOWNTO 0);
	sub_wire8    <= data10x(0 DOWNTO 0);
	sub_wire7    <= data11x(0 DOWNTO 0);
	sub_wire6    <= data12x(0 DOWNTO 0);
	sub_wire5    <= data13x(0 DOWNTO 0);
	sub_wire4    <= data14x(0 DOWNTO 0);
	sub_wire3    <= data15x(0 DOWNTO 0);
	result    <= sub_wire0(5 DOWNTO 0);
	sub_wire1    <= data16x(0 DOWNTO 0);
	sub_wire2(16, 0)    <= sub_wire1(0);
	sub_wire2(15, 0)    <= sub_wire3(0);
	sub_wire2(14, 0)    <= sub_wire4(0);
	sub_wire2(13, 0)    <= sub_wire5(0);
	sub_wire2(12, 0)    <= sub_wire6(0);
	sub_wire2(11, 0)    <= sub_wire7(0);
	sub_wire2(10, 0)    <= sub_wire8(0);
	sub_wire2(9, 0)    <= sub_wire9(0);
	sub_wire2(8, 0)    <= sub_wire10(0);
	sub_wire2(7, 0)    <= sub_wire11(0);
	sub_wire2(6, 0)    <= sub_wire12(0);
	sub_wire2(5, 0)    <= sub_wire13(0);
	sub_wire2(4, 0)    <= sub_wire14(0);
	sub_wire2(3, 0)    <= sub_wire15(0);
	sub_wire2(2, 0)    <= sub_wire16(0);
	sub_wire2(1, 0)    <= sub_wire17(0);
	sub_wire2(0, 0)    <= sub_wire18(0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 0,
		representation => "UNSIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 17,
		width => 1,
		widthr => 6,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "17"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "6"
-- Retrieval info: USED_PORT: data0x 0 0 1 0 INPUT NODEFVAL "data0x[0..0]"
-- Retrieval info: USED_PORT: data10x 0 0 1 0 INPUT NODEFVAL "data10x[0..0]"
-- Retrieval info: USED_PORT: data11x 0 0 1 0 INPUT NODEFVAL "data11x[0..0]"
-- Retrieval info: USED_PORT: data12x 0 0 1 0 INPUT NODEFVAL "data12x[0..0]"
-- Retrieval info: USED_PORT: data13x 0 0 1 0 INPUT NODEFVAL "data13x[0..0]"
-- Retrieval info: USED_PORT: data14x 0 0 1 0 INPUT NODEFVAL "data14x[0..0]"
-- Retrieval info: USED_PORT: data15x 0 0 1 0 INPUT NODEFVAL "data15x[0..0]"
-- Retrieval info: USED_PORT: data16x 0 0 1 0 INPUT NODEFVAL "data16x[0..0]"
-- Retrieval info: USED_PORT: data1x 0 0 1 0 INPUT NODEFVAL "data1x[0..0]"
-- Retrieval info: USED_PORT: data2x 0 0 1 0 INPUT NODEFVAL "data2x[0..0]"
-- Retrieval info: USED_PORT: data3x 0 0 1 0 INPUT NODEFVAL "data3x[0..0]"
-- Retrieval info: USED_PORT: data4x 0 0 1 0 INPUT NODEFVAL "data4x[0..0]"
-- Retrieval info: USED_PORT: data5x 0 0 1 0 INPUT NODEFVAL "data5x[0..0]"
-- Retrieval info: USED_PORT: data6x 0 0 1 0 INPUT NODEFVAL "data6x[0..0]"
-- Retrieval info: USED_PORT: data7x 0 0 1 0 INPUT NODEFVAL "data7x[0..0]"
-- Retrieval info: USED_PORT: data8x 0 0 1 0 INPUT NODEFVAL "data8x[0..0]"
-- Retrieval info: USED_PORT: data9x 0 0 1 0 INPUT NODEFVAL "data9x[0..0]"
-- Retrieval info: USED_PORT: result 0 0 6 0 OUTPUT NODEFVAL "result[5..0]"
-- Retrieval info: CONNECT: @data 1 0 1 0 data0x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 10 1 0 data10x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 11 1 0 data11x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 12 1 0 data12x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 13 1 0 data13x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 14 1 0 data14x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 15 1 0 data15x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 16 1 0 data16x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 1 1 0 data1x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 2 1 0 data2x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 3 1 0 data3x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 4 1 0 data4x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 5 1 0 data5x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 6 1 0 data6x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 7 1 0 data7x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 8 1 0 data8x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 9 1 0 data9x 0 0 1 0
-- Retrieval info: CONNECT: result 0 0 6 0 @result 0 0 6 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_parallelAdder.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_parallelAdder.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_parallelAdder.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_parallelAdder.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_parallelAdder_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf

library verilog;
use verilog.vl_types.all;
entity Arena_register_vlg_vec_tst is
end Arena_register_vlg_vec_tst;

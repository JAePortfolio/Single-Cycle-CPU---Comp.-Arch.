library verilog;
use verilog.vl_types.all;
entity Arena_32bit_divider_usingVHDL_vlg_vec_tst is
end Arena_32bit_divider_usingVHDL_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_3to8Decoder_vlg_vec_tst is
end Arena_3to8Decoder_vlg_vec_tst;

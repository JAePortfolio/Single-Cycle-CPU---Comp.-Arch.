library verilog;
use verilog.vl_types.all;
entity Arena_Control_vlg_vec_tst is
end Arena_Control_vlg_vec_tst;

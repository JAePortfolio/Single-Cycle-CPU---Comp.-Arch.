library verilog;
use verilog.vl_types.all;
entity Arena_8to3Encoder_vlg_vec_tst is
end Arena_8to3Encoder_vlg_vec_tst;

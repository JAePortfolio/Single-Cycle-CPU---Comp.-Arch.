library verilog;
use verilog.vl_types.all;
entity Arena_HalfAdder_vlg_vec_tst is
end Arena_HalfAdder_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_32bitAccumulator_withSegmentDisplay_vlg_check_tst is
    port(
        AccumOut        : in     vl_logic_vector(31 downto 0);
        Arena_A         : in     vl_logic_vector(31 downto 0);
        Arena_AccumOut_32bit: in     vl_logic_vector(31 downto 0);
        Arena_Bout_32bit: in     vl_logic;
        Arena_Cout_32bit: in     vl_logic;
        Arena_segment1_A: in     vl_logic;
        Arena_segment1_B: in     vl_logic;
        Arena_segment1_C: in     vl_logic;
        Arena_segment1_D: in     vl_logic;
        Arena_segment1_E: in     vl_logic;
        Arena_segment1_F: in     vl_logic;
        Arena_segment1_G: in     vl_logic;
        Arena_segment2_A: in     vl_logic;
        Arena_segment2_B: in     vl_logic;
        Arena_segment2_C: in     vl_logic;
        Arena_segment2_D: in     vl_logic;
        Arena_segment2_E: in     vl_logic;
        Arena_segment2_F: in     vl_logic;
        Arena_segment2_G: in     vl_logic;
        Arena_segment3_A: in     vl_logic;
        Arena_segment3_B: in     vl_logic;
        Arena_segment3_C: in     vl_logic;
        Arena_segment3_D: in     vl_logic;
        Arena_segment3_E: in     vl_logic;
        Arena_segment3_F: in     vl_logic;
        Arena_segment3_G: in     vl_logic;
        Arena_segment4_A: in     vl_logic;
        Arena_segment4_B: in     vl_logic;
        Arena_segment4_C: in     vl_logic;
        Arena_segment4_D: in     vl_logic;
        Arena_segment4_E: in     vl_logic;
        Arena_segment4_F: in     vl_logic;
        Arena_segment4_G: in     vl_logic;
        Arena_segment5_A: in     vl_logic;
        Arena_segment5_B: in     vl_logic;
        Arena_segment5_C: in     vl_logic;
        Arena_segment5_D: in     vl_logic;
        Arena_segment5_E: in     vl_logic;
        Arena_segment5_F: in     vl_logic;
        Arena_segment5_G: in     vl_logic;
        Arena_segment6_A: in     vl_logic;
        Arena_segment6_B: in     vl_logic;
        Arena_segment6_C: in     vl_logic;
        Arena_segment6_D: in     vl_logic;
        Arena_segment6_E: in     vl_logic;
        Arena_segment6_F: in     vl_logic;
        Arena_segment6_G: in     vl_logic;
        Arena_segment7_A: in     vl_logic;
        Arena_segment7_B: in     vl_logic;
        Arena_segment7_C: in     vl_logic;
        Arena_segment7_D: in     vl_logic;
        Arena_segment7_E: in     vl_logic;
        Arena_segment7_F: in     vl_logic;
        Arena_segment7_G: in     vl_logic;
        Arena_segment8_A: in     vl_logic;
        Arena_segment8_B: in     vl_logic;
        Arena_segment8_C: in     vl_logic;
        Arena_segment8_D: in     vl_logic;
        Arena_segment8_E: in     vl_logic;
        Arena_segment8_F: in     vl_logic;
        Arena_segment8_G: in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_32bitAccumulator_withSegmentDisplay_vlg_check_tst;

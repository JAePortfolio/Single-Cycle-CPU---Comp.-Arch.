library verilog;
use verilog.vl_types.all;
entity Arena_16bitMultiplier_withSegmentDisplay_vlg_vec_tst is
end Arena_16bitMultiplier_withSegmentDisplay_vlg_vec_tst;

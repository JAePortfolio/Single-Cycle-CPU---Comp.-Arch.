library verilog;
use verilog.vl_types.all;
entity Arena_bitwise_setLessThanUnsigned_vlg_check_tst is
    port(
        Arena_result_sltuOUT: in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_bitwise_setLessThanUnsigned_vlg_check_tst;

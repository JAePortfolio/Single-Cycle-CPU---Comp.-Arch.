library verilog;
use verilog.vl_types.all;
entity Arena_SRAM_vlg_vec_tst is
end Arena_SRAM_vlg_vec_tst;

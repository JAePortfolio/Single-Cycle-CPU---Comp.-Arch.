library verilog;
use verilog.vl_types.all;
entity Arena_bitwise_setLessThanSigned_vlg_vec_tst is
end Arena_bitwise_setLessThanSigned_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_1bitDivider_vlg_vec_tst is
end Arena_1bitDivider_vlg_vec_tst;

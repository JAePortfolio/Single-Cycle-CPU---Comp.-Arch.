library verilog;
use verilog.vl_types.all;
entity Arena_fullSubtractor_vlg_vec_tst is
end Arena_fullSubtractor_vlg_vec_tst;

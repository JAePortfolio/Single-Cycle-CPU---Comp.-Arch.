library verilog;
use verilog.vl_types.all;
entity Arena_bitwiseand_vlg_vec_tst is
end Arena_bitwiseand_vlg_vec_tst;

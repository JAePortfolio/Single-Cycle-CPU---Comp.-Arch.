library verilog;
use verilog.vl_types.all;
entity Arena_Sign_Extend_16to32_vlg_vec_tst is
end Arena_Sign_Extend_16to32_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_16bitFullAdder_vlg_vec_tst is
end Arena_16bitFullAdder_vlg_vec_tst;

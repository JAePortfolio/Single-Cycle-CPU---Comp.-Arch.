library verilog;
use verilog.vl_types.all;
entity Arena_simpleCircuit_vlg_vec_tst is
end Arena_simpleCircuit_vlg_vec_tst;

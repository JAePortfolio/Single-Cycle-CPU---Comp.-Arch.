library verilog;
use verilog.vl_types.all;
entity Arena_4to16Decoder_vlg_vec_tst is
end Arena_4to16Decoder_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_bitwisexor_vlg_vec_tst is
end Arena_bitwisexor_vlg_vec_tst;

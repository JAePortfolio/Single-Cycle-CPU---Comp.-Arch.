library verilog;
use verilog.vl_types.all;
entity Arena_bitwiseOperation_decoder_vlg_vec_tst is
end Arena_bitwiseOperation_decoder_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_mux2to1_vlg_vec_tst is
end Arena_mux2to1_vlg_vec_tst;

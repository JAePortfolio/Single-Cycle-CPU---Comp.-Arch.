library verilog;
use verilog.vl_types.all;
entity Single_Cycle_CPU_withDisplays_vlg_vec_tst is
end Single_Cycle_CPU_withDisplays_vlg_vec_tst;

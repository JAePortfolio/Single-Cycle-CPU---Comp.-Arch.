library verilog;
use verilog.vl_types.all;
entity Arena_bitrotationleft_vlg_vec_tst is
end Arena_bitrotationleft_vlg_vec_tst;

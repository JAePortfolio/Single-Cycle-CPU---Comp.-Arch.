library verilog;
use verilog.vl_types.all;
entity Arena_SRAM_vlg_check_tst is
    port(
        Arena_OUT       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_SRAM_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_bitwisenot_vlg_vec_tst is
end Arena_bitwisenot_vlg_vec_tst;

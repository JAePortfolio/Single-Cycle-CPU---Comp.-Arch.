library verilog;
use verilog.vl_types.all;
entity Arena_16x32_SRAM_vlg_vec_tst is
end Arena_16x32_SRAM_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_DLatch_vlg_vec_tst is
end Arena_DLatch_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_4bit_arrayMultipler_vlg_vec_tst is
end Arena_4bit_arrayMultipler_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_D_FlipFlop_vlg_vec_tst is
end Arena_D_FlipFlop_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_ProgramCounter_32bit_vlg_vec_tst is
end Arena_ProgramCounter_32bit_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_16bitMultiplier_using_registers_v1_vlg_vec_tst is
end Arena_16bitMultiplier_using_registers_v1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_mux2to1_vlg_check_tst is
    port(
        Arena_M         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_mux2to1_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_simpleCircuit_vlg_check_tst is
    port(
        Arena_F         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_simpleCircuit_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_bitshiftleft_vlg_vec_tst is
end Arena_bitshiftleft_vlg_vec_tst;

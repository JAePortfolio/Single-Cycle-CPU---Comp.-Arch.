library verilog;
use verilog.vl_types.all;
entity Arena_bitshiftright_vlg_vec_tst is
end Arena_bitshiftright_vlg_vec_tst;

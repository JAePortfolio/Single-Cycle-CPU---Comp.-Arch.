-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: Arena_muxLPM.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY Arena_muxLPM IS
	PORT
	(
		Arena_data0		: IN STD_LOGIC ;
		Arena_data1		: IN STD_LOGIC ;
		Arena_sel		: IN STD_LOGIC ;
		Arena_result		: OUT STD_LOGIC 
	);
END Arena_muxLPM;


ARCHITECTURE SYN OF arena_muxlpm IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL Arena_sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL Arena_sub_wire1	: STD_LOGIC ;
	SIGNAL Arena_sub_wire2	: STD_LOGIC ;
	SIGNAL Arena_sub_wire3	: STD_LOGIC_2D (1 DOWNTO 0, 0 DOWNTO 0);
	SIGNAL Arena_sub_wire4	: STD_LOGIC ;
	SIGNAL Arena_sub_wire5	: STD_LOGIC ;
	SIGNAL Arena_sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);

BEGIN
	Arena_sub_wire4    <= Arena_data0;
	Arena_sub_wire1    <= Arena_sub_wire0(0);
	Arena_result    <= Arena_sub_wire1;
	Arena_sub_wire2    <= Arena_data1;
	Arena_sub_wire3(1, 0)    <= Arena_sub_wire2;
	Arena_sub_wire3(0, 0)    <= Arena_sub_wire4;
	Arena_sub_wire5    <= Arena_sel;
	Arena_sub_wire6(0)    <= Arena_sub_wire5;

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 2,
		lpm_type => "LPM_MUX",
		lpm_width => 1,
		lpm_widths => 1
	)
	PORT MAP (
		data => Arena_sub_wire3,
		sel => Arena_sub_wire6,
		result => Arena_sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
-- Retrieval info: USED_PORT: data0 0 0 0 0 INPUT NODEFVAL "data0"
-- Retrieval info: USED_PORT: data1 0 0 0 0 INPUT NODEFVAL "data1"
-- Retrieval info: USED_PORT: result 0 0 0 0 OUTPUT NODEFVAL "result"
-- Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL "sel"
-- Retrieval info: CONNECT: @data 1 0 1 0 data0 0 0 0 0
-- Retrieval info: CONNECT: @data 1 1 1 0 data1 0 0 0 0
-- Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 0 0 @result 0 0 1 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_muxLPM.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_muxLPM.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_muxLPM.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_muxLPM.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Arena_muxLPM_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm

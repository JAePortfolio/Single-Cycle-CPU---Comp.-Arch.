library verilog;
use verilog.vl_types.all;
entity Arena_FullAdder_vlg_vec_tst is
end Arena_FullAdder_vlg_vec_tst;

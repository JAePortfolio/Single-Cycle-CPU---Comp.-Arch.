library verilog;
use verilog.vl_types.all;
entity Arena_32bitInput_vlg_vec_tst is
end Arena_32bitInput_vlg_vec_tst;

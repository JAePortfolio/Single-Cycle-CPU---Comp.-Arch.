library verilog;
use verilog.vl_types.all;
entity Arena_muxLPM_vlg_vec_tst is
end Arena_muxLPM_vlg_vec_tst;

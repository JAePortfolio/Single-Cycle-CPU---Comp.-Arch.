library verilog;
use verilog.vl_types.all;
entity Arena_D_FlipFlop_vlg_check_tst is
    port(
        Arena_Q         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Arena_D_FlipFlop_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Arena_SRLatch_vlg_vec_tst is
end Arena_SRLatch_vlg_vec_tst;

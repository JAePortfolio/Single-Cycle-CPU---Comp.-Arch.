library verilog;
use verilog.vl_types.all;
entity Arena_bitrotationright_vlg_vec_tst is
end Arena_bitrotationright_vlg_vec_tst;
